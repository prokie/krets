
V1 in_ac1 0 SIN(0 5 60 0 0 0)
V2 in_ac2 0 SIN(0 -5 60 0 0 0)

D1 in_ac1 out_dc DMOD
D2 in_ac2 out_dc DMOD  
D3 0 in_ac1 DMOD
D4 0 in_ac2 DMOD

C1 out_dc 0 100u
R1 out_dc 0 1k 

.model DMOD D (is=1e-12)

.control
  tran 0.1ms 50ms
  run
  plot v(in_ac1,in_ac2) v(out_dc)
.endc
.end