* Simple diode circuit for DC analysis
V1 in 0 1
R1 in out 1000
D1 out 0 DMOD


.model DMOD D



.control
options abstol=1e-12 reltol=1e-6
dc V1 0 2.0 0.01
save all
print all
.endc

